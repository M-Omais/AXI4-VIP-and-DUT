package tx_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "tx_item.sv"
    `include "axi_seqs.sv"
    `include "axi_sequencer.sv"
    `include "axi_driver.sv"
    `include "axi_monitor.sv"
    `include "axi_agent.sv"
    `include "axi_sb.sv"
    `include "axi_env.sv"
    `include "Test.sv"
endpackage