package seq_pkg;
	import uvm_pkg::*;
    `include "uvm_macros.svh"
	`include "tx_item.sv"
    `include "write_seq.sv"
    `include "read_seq.sv"
    `include "fixed_burst.sv"
    `include "incr_burst.sv"
    `include "warp_burst.sv"
endpackage
